library IEEE;
use IEEE.Std_Logic_1164.all;
use IEEE.std_logic_signed.all; -- Para poder usar o operador +

entity topo is
port(CLOCK_50:in std_logic;
     CLK_500Hz:in std_logic;
     KEY:in std_logic_vector(3 downto 0);
     SW:in std_logic_vector(17 downto 0);
     LEDR:out std_logic_vector(17 downto 0);
     HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7: out std_logic_vector(6 downto 0));
end topo;

architecture circuito_exe2 of topo is
signal A, F, F1, F2, F3, F4: std_logic_vector(3 downto 0); --vetores intermediários
signal C: std_logic_vector(1 downto 0); --vetores intermediários

component mux4_1 is
port (F1,F2,F3,F4: in std_logic_vector(3 downto 0);
sel: in std_logic_vector(1 downto 0);
F: out std_logic_vector(3 downto 0)
);
end component;

component mux2_1 is
port (
F1: in std_logic_vector(6 downto 0);
F2: in std_logic_vector(6 downto 0);
sel: in std_logic;
F: out std_logic_vector(6 downto 0)
);
end component;

component decod_C2 is
port (G: in std_logic_vector(3 downto 0);
F: out std_logic_vector(6 downto 0)
);
end component;

component  decod is
port (C: in std_logic_vector(1 downto 0);
F: out std_logic_vector(6 downto 0)
);
end component;

begin

A <= SW(3 downto 0);
C <= SW(9 downto 8);

MUX4: mux4_1 port map((A+4),(A+5), (A-2), (A-1), SW(9 downto 8), F);

MUX2a: mux2_1 port map("1111111", "0111111", SW(3), HEX6);
MUX2b: mux2_1 port map("0001111", "0111111", SW(9), HEX4);
MUX2c: mux2_1 port map("1111111", "0111111", F(3), HEX1);

DEC2a: decod_C2 port map(SW(3 downto 0), HEX5);
DEC2b: decod_C2 port map(F, HEX0);

DEC: decod port map(SW(9 downto 8), HEX3);

HEX2 <= "0110111";

end circuito_exe2;
